`ifndef IMMCODE
`define IMMCODE

`define IMM_R_TYPE 3'b000
`define IMM_I_TYPE 3'b001
`define IMM_S_TYPE 3'b010
`define IMM_B_TYPE 3'b011
`define IMM_U_TYPE 3'b100
`define IMM_JAL    3'b101
`define IMM_JALR   3'b110
`define IMM_CSR    3'b111

`endif //IMMCODE
