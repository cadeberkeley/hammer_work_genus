/bwrcq/scratch/caderichard/hammer/hammer/technology/asap7/sram_compiler/memories/lef/SRAM2RW32x8_x4.lef