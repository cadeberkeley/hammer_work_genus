`ifndef LOADOP
`define LOADOP

`define FUNCT3_LB	3'b000
`define FUNCT3_LH	3'b001
`define FUNCT3_LW	3'b010
`define FUNCT3_LBU	3'b100
`define FUNCT3_LHU	3'b101
`define FUNCT3_LWU	3'b110

`define SEL_LW	2'b00
`define SEL_LH	2'b01
`define SEL_LB	2'b10

`endif //LOADOP
