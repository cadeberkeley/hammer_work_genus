`ifndef STOREOP
`define STOREOP

`define FUNCT3_SW	3'b010
`define FUNCT3_SH	3'b001
`define FUNCT3_SB	3'b000

`endif // STOREOP
