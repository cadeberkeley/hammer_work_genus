/bwrcq/B/asap7/asap7sc7p5t_27/techlef_misc/asap7_tech_4x_201209.lef