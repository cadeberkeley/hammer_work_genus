/bwrcq/scratch/caderichard/hammer/hammer/technology/asap7/sram_compiler/memories/lef/SRAM1RW4096x16_x4.lef